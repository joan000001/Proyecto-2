module keypad_scan #(
    
)(
    input  logic        clk,
    input  logic        rst_n,
    input  logic [3:0]  columnas,
    output logic [3:0]  filas,
    output logic [1:0]  row,
    output logic [1:0]  col,
    output logic        valid
);



endmodule