module top (
    input  logic        clk,
    input  logic [3:0]  columnas,
    output logic [3:0]  filas,
    output logic [6:0]  segments,
    output logic [2:0]  enable_displays
);


endmodule